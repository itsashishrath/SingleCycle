module Mux(
	input [31:0]SignImm,
	input [31:] A3,
	input sel)