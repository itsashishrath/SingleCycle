module regFile(
	input clk,
	input A1,
	input A2,
	input A3
	input WD3,
	input WE3,
	output RD2,