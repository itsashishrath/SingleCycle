module PC(
	input clk,
	output[31:0] pc_out,
	input [31:0] pc_in);

	reg [31:0] instr_temp=instr_in;
	

	


	