module InstrMem(
	input [31:0]A,
	output [31:0] RD
	);
	
	reg [15:0]PC
	
//	address A usjagah se 32 bit ka instruction lena 
	
//	RD=instruction;
	
